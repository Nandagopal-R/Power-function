`timescale 1ns / 1ps
module pow2(ip,out,clk);
reg [31:0] a [12:0],b [12:0],c[11:0];
reg [31:0] z;
wire [31:0] y;
reg [31:0] exp;  //,ip=32'b00111111000100010110100001110011;   //0.568
input [31:0] ip;
output reg [31:0] out;
input clk;

wire [31:0] op1,op2,op3,op4,op5,op;
reg[3:0] i=0,j;
reg [2:0] k=0,l=0,m=0;

always@(posedge clk)
begin

a[0]=32'b00000000000000000000000000000000;    //0
a[1]=32'b00111110000000000000000000000000;    //0.125
a[2]=32'b00111110011100000000011010001110;    //0.2344
a[3]=32'b00111110101010010000001011011110;    //0.3301
a[4]=32'b00111110110100111101110110011000;    //0.4138
a[5]=32'b00111110111110010110010100101100;    //0.4871
a[6]=32'b00111111000011010001101101110001;    //0.5512;
a[7]=32'b00111111000110110111100000000011;    //0.6073;
a[8]=32'b00111111001101001001101110100110;    //0.7055;
a[9]=32'b00111111010001110111001100011001;    //0.7791;
a[10]=32'b00111111010101011001010010101111;   //0.8343;
a[11]=32'b00111111011010101100110110011111;   //0.9172;
a[12]=32'b00111111100000000000000000000000;   //1;

 

b[0]=32'b00111111100000000000000000000000;   //1
b[1]=32'b00111111100010111001010110111100;   //1.090507
b[2]=32'b00111111100101101001010011010101;   //1.176417
b[3]=32'b00111111101000001110100010100111;   //1.257100
b[4]=32'b00111111101010101000010100110100;   //1.332190;
b[5]=32'b00111111101100110110100001101010;   //1.401624;
b[6]=32'b00111111101110111000111100001100;   //1.465303;
b[7]=32'b00111111110000101111111011101111;   //1.523405;
b[8]=32'b00111111110100001011101100010011;   //1.630709;
b[9]=32'b00111111110110111010011111011011;   //1.716060;
b[10]=32'b00111111111001000011100100001101;  //1.782991;
b[11]=32'b00111111111100011011100010011001;  //1.888446;
b[12]=32'b01000000000000000000000000000000;  //2.0;



c[0]=32'b01000001000000000000000000000000;    //8
c[1]=32'b01000001000100100100000001001111;    //9.1407
c[2]=32'b01000001001001110011000001010101;    //10.4493
c[3]=32'b01000001001111110010100010001101;    //11.9474
c[4]=32'b01000001010110100100011110101110;    //13.6425
c[5]=32'b01000001011110011001110000001111;    //15.6006
c[6]=32'b01000001100011101001101000110111;    //17.8253
c[7]=32'b01000001001000101110111001100011;    //10.1832
c[8]=32'b01000001010110010110001111110001;    //13.5869;
c[9]=32'b01000001100100001110110101011101;    //18.1159;
c[10]=32'b01000001010000010000000011010010;   //12.0627;
c[11]=32'b01000001010000010011110000110110;   //12.0772;


for(i=0;i<12;i=i+1)
begin
if(ip>=a[i] && ip<=a[i+1])
begin
j=i;
end
end
out=in5.c;
end

subt in1(b[j],b[j+1],op1);
mul in2(op1,c[j],op2);
subt in3(a[j],ip,op3);
mul in4(op2,op3,op4);
add in5(op4,b[j],op);

endmodule







