`timescale 1ns / 1ps
module log2(user_ip,out,clk);
reg [31:0] a [13:0],b [13:0],c[13:0];
reg [31:0] z;
wire [31:0] y;
output reg [31:0] out;

reg [31:0] ip;   
input [31:0] user_ip;                           
reg [32:0] cnst=32'b01000010111111100000000000000000;
reg [31:0] exp;
input clk;
wire [31:0] op1,op2,op3,op4,op5,op;
integer i,j,k,l,m;

always@(posedge clk)
begin
a[0]= 32'b00111111100000000000000000000000;    //1
a[1]= 32'b00111111100010000000000000000000;    //1.0625
a[2]= 32'b00111111100011111000000000110100;    //1.1211
a[3]= 32'b00111111100101101000011100101011;    //1.1760
a[4]= 32'b00111111100111010001111010111000;    //1.2275
a[5]= 32'b00111111101000110100110101101010;    //1.2758
a[6]= 32'b00111111101011101000000010011101;    //1.3663;
a[7]= 32'b00111111101110010000011000100101;    //1.4455;
a[8]= 32'b00111111110000011110010011110111;    //1.5148;
a[9]= 32'b00111111110010011010100111111100;    //1.5755;
a[10]=32'b00111111110101110011111010101011;   //1.6816;
a[11]=32'b00111111111000010110111100000000;   //1.7612;
a[12]=32'b00111111111100001011011110000000;   //1.8806;
a[13]=32'b01000000000000000000000000000000;   //2;

b[0]= 32'b00000000000000000000000000000000;   //0
b[1]= 32'b00111101101100110011001100110011;   //0.0875
b[2]= 32'b00111110001010001101101110001100;   //0.1649
b[3]= 32'b00111110011011111000001101111011;   //0.2339
b[4]= 32'b00111110100101110111001100011001;   //0.2958;
b[5]= 32'b00111110101100111110101010110011;   //0.3514;
b[6]= 32'b00111110111001101000110110111001;   //0.4503;
b[7]= 32'b00111111000010000001011011110000;   //0.5316;
b[8]= 32'b00111111000110010110010100101100;   //0.5992;
b[9]= 32'b00111111001001111110001010000010;   //0.6558;
b[10]=32'b00111111001111111111001011100101;  //0.7498;
b[11]=32'b00111111010100010000110010110011;  //0.8166;
b[12]=32'b00111111011010010100010001100111;  //0.9112;
b[13]=32'b00111111100000000000000000000000;  //1;

c[0]= 32'b00111111110011001100110011001101;    //1.6
c[1]= 32'b01000001100010001000010010110110;    //17.0648
c[2]= 32'b01000001100100011011100000011101;    //18.2149
c[3]= 32'b01000001100110110101011011010110;    //19.4174
c[4]= 32'b01000001101001011010000110101000;    //20.7039;
c[5]= 32'b01000001001100001100101110101010;    //11.0497;
c[6]= 32'b01000001010010100000010100101100;    //12.6262;
c[7]= 32'b01000001011001101110000101010111;    //14.4300;
c[8]= 32'b01000001100000111100101110110100;    //16.4744;
c[9]= 32'b01000001000101101100110100010111;    //9.4250;
c[10]=32'b01000001010010010000000101001001;   //12.5628;
c[11]=32'b01000001000001100000000011011011;   //8.3752;
c[12]=32'b01000001000011000101100111010011;   //8.77192
c[13]=32'b00111111100000000000000000000000;   //1;

ip[31]=0;
ip[30:23]=8'b01111111;
ip[22:0]=user_ip[22:0];

exp[31]=0;


for(l=0;l<8;l=l+1)
begin
if(user_ip[23+l]==1)
k=l;
end

if(k==7)
begin
exp[30:23]=8'b10000110;
exp[22:16]=user_ip[29:23];
exp[15:0]=0;
end

if(k==6)
begin
exp[30:23]=8'b10000101;
exp[22:17]=user_ip[28:23];
exp[16:0]=0;
end

if(k==5)
begin
exp[30:23]=8'b10000100;
exp[22:18]=user_ip[27:23];
exp[17:0]=0;
end

if(k==4)
begin
exp[30:23]=8'b10000011;
exp[22:19]=user_ip[26:23];
exp[18:0]=0;
end

if(k==3)
begin
exp[30:23]=8'b10000010;
exp[22:20]=user_ip[25:23];
exp[19:0]=0;
end

if(k==2)
begin
exp[30:23]=8'b10000001;
exp[22:21]=user_ip[24:23];
exp[20:0]=0;
end


/*
ip[0]=32'b00111111100100110011001100110011;    //1.15-correct
ip[1]=32'b00111111101000010100011110101110;    //1.26-correct
ip[2]=32'b00111111111100000010000011000101;     //1.876-correct
ip[3]=32'b00111111111101101010011111110000;     //1.927
*/

for(i=0;i<13;i=i+1)
begin
if(ip>=a[i] && ip<=a[i+1])
begin

j=i;
end
end
out=in7.c;
//w=w+1;
end



//conv in0(user_ip,ip,exp,clk);
subt in1(b[j],b[j+1],op1,clk);
mul in2(op1,c[j],op2,clk);
subt in3(a[j],ip,op3,clk);
mul in4(op2,op3,op4,clk);
add in5(op4,b[j],op,clk);
subt in6(cnst,exp,op5,clk);
add in7(op,op5,y,clk);


endmodule







